`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    13:12:10 04/03/2023 
// Design Name: 
// Module Name:    ZMux10to1 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module ZPulseCounter_Mux10to1(
    input clk,
    input rst_n,
    input [3:0] select,
    output [3:0] dout
    );


endmodule
