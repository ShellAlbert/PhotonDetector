`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    08:39:26 03/20/2023 
// Design Name: 
// Module Name:    ZOLED_Module_MapY2Page 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module ZOLED_Module_MapY2Page(
    input clk,
    input rst_n,
    input iY,
    output [7:0] oPage,
    output [7:0] oBitMask
    );


endmodule
