`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    13:38:26 02/22/2023 
// Design Name: 
// Module Name:    ZKey_Module_Delay 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module ZKey_Module_Delay(
    input clk,
    input rst_n,
    input en,
    input pulse,
    output delayed_pulse
    );


endmodule
