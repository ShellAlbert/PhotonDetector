`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    10:44:26 02/22/2023 
// Design Name: 
// Module Name:    ZKey_Module_Edge_Detector 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module ZKey_Module_Edge_Detector(
    input clk,
    input rst_n,
    input key_pin,
    output h2l_edge,
    output l2h_edge
    );


endmodule
