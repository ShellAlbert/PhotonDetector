`timescale 10ns/1ns
module ZPhotonDetector_tb;

reg iPulse;
reg iSync50Hz;

initial begin
    
end

endmodule
