`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    14:28:58 04/25/2023 
// Design Name: 
// Module Name:    zpush_button 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module zpush_button(
    input clk,
    input rst_n,
    input en,
    input [3:0] iButton,
    output [3:0] oButton
    );


endmodule
