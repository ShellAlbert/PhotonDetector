`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    09:15:57 04/20/2023 
// Design Name: 
// Module Name:    ZShift_and_Draw 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
`include "../ColorTable/ZRGB565_ColorTable.v"
module ZShift_and_Draw(
    input clk,
    input rst_n,
    input en,

	//New PulseCounter comes.
	input iDataUpdate,
	input [15:0] iPulseCounter,
    
	//SDRAM Read Glue Logic.
    output reg [23:0] oSDRAM_Rd_Addr, //output, Bank(2)+Row(13)+Column(9)=(24)
    input [15:0] iSDRAM_Data, //input, read back data from SDRAM.

    output reg oSDRAM_Rd_Req, //output, [1]=1:Write, [0]=1:Read.
    input iSDRAM_Rd_Done, //input,[1]=1:write done, [0]=1:read done.

	//SDRAM Write Glue Logic.
    output reg [23:0] oSDRAM_Wr_Addr, //output, Bank(2)+Row(13)+Column(9)=(24)
    output reg [15:0] oSDRAM_Wr_Data, //ouptut, write data to SDRAM.

    output reg oSDRAM_Wr_Req, //output, [1]=1:Write, [0]=1:Read.
    input iSDRAM_Wr_Done //input, SDRAM write done signal.
    );

//SDRAM Space Assignment
//0~383999: (480*800-1): LCD GRAM. 
//384000~384599: (384000+600-1): Photon Counter.

//Lock in new pulse counter.
reg [15:0] lockInPulseCounter;
always @(posedge clk or negedge rst_n)
if(!rst_n)	begin
				lockInPulseCounter<=0;
			end
else if(iDataUpdate)	begin
							lockInPulseCounter<=iPulseCounter;
						end
//Do shift movement.
//Eliminate the oldest value and add the new pulse counter.
//Left Shift Effect.
reg [31:0] i;
reg [31:0] ringbuffer_wr_addr;
reg [15:0] CNT1;
reg [31:0] ringbuffer_rd_addr;

reg [15:0] newPulseCounter;
reg [31:0] GRAM_X;
reg [31:0] GRAM_Y;
reg [15:0] CNT2;
always @(posedge clk or negedge rst_n)
if(!rst_n)	begin
				i<=0;
				CNT1<=0;
				CNT2<=0;
				
				//SDRAM Read.
				oSDRAM_Rd_Req<=0;
				oSDRAM_Rd_Addr<=0;

				//SDRAM Write.
				oSDRAM_Wr_Req<=0;
				oSDRAM_Wr_Addr<=0;
				oSDRAM_Wr_Data<=0;

				newPulseCounter<=0;
				ringbuffer_wr_addr<=384000;
			end
else if(en) begin
			case(i)
				0: //Write the new pulse counter to 384600.
				//384000,384000+1,384000+2,384000+3, ... ... 384000+599,384000+600.
				//Left Shift the entire area, so we should write the new pulse couter to 384000+600.
				//Ring buffer to write new pulse counter to SDRAM.
					if(iSDRAM_Wr_Done) begin 
											oSDRAM_Wr_Req<=0; 
											i<=i+1'b1; 
										end
					else begin 
							oSDRAM_Wr_Req<=1; 
							oSDRAM_Wr_Addr<=ringbuffer_wr_addr;
							oSDRAM_Wr_Data<=iPulseCounter;
						end
				1: //Ring buffer to loop.
					begin
						if(ringbuffer_wr_addr==384599) 
							ringbuffer_wr_addr<=384000; 
						else 
							ringbuffer_wr_addr<=ringbuffer_wr_addr+1'b1; 
						/////////////////
						i<=i+1'b1;
					end
				2: //read from ring buffer and write GRAM.
					if(1/*newPulseCounter!=lockInPulseCounter*/) begin
															ringbuffer_rd_addr<=384000;
															
															//GRAM Plain yOffset=20*480=9600.
															GRAM_Y<=9600;
															i<=i+1'b1;
														end
				3: //Read from ring buffer.
					if(iSDRAM_Rd_Done) begin 
										oSDRAM_Rd_Req<=1'b0; 
										//GRAM X.
										GRAM_X<=10+iSDRAM_Data>>1; //+xOffset.
										CNT1<=iSDRAM_Data>>1;//iSDRAM_Data;
										i<=i+1'b1; 
									end
					else begin 
							oSDRAM_Rd_Req<=1'b1; 
							oSDRAM_Rd_Addr<=ringbuffer_rd_addr;
						end
				4: //GRAM: Write to GRAM the toppest point.
					if(iSDRAM_Wr_Done) begin 
											oSDRAM_Wr_Req<=0; 
											i<=i+1'b1; 
										end
					else begin 
							oSDRAM_Wr_Req<=1;
							oSDRAM_Wr_Addr<=GRAM_Y+GRAM_X-1;
							oSDRAM_Wr_Data<=`Color_Pink;
						end
				5: //GRAM: Loop to draw from top to bottom to generate histogram.
					if(CNT1==0) begin i<=i+1'b1; end
					else begin 
							CNT1<=CNT1-1'b1; 
							GRAM_X<=GRAM_X-1'b1; 
							i<=i-1'b1; 
						end
				6: //Loop 600-1=599 times.
					if(CNT2==599) begin CNT2<=0; i<=i+1'b1; end
					else begin 
							CNT2<=CNT2+1'b1; 
							ringbuffer_rd_addr<=ringbuffer_rd_addr+1'b1;
							//GRAM Y. Next Y.
							GRAM_Y<=GRAM_Y+480; 
							i<=3; //Loop to write GRAM.
						end
				7: //
					begin i<=0; end
			endcase
		 end
endmodule
