`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    11:04:46 04/02/2023 
// Design Name: 
// Module Name:    ZRTC_Counter 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module ZRTC_Counter(
    input clk,
    input rst_n,
    input en,
    output [5:0] hour,
    output [5:0] minute,
    output [5:0] second
    );


endmodule
