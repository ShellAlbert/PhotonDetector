`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 10/24/2023 10:46:31 AM
// Design Name: 
// Module Name: ZPower_EN
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module ZPower_EN(
    input iClk,
    input iRst_N,
    output oEn
    );
assign oEn=1'b1;
endmodule
