`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    13:48:41 04/06/2023 
// Design Name: 
// Module Name:    ZExSignalSync 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module ZExSignalSync(
    input clk,
    input rst_n,
    input sig_in,
    output sig_out
    );


endmodule
