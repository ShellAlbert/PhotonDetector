`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    11:05:09 10/29/2022 
// Design Name: 
// Module Name:    ZsyDotMatrix 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module ZsyDotMatrix(
    input clk,
    input rst_n,
    input [4:0] addr,
    output [127:0] data_top,
	output [127:0] data_btm
    );

reg [127:0] rdata_top;
reg [127:0] rdata_btm;
always @ (posedge clk or negedge rst_n)
if(!rst_n)	begin
				rdata_top<=128'd0;
				rdata_btm<=128'd0;
			end
else case(addr)
		5'd0:begin
//{00_00_F8_49_4A_4C_48_F8_48_4C_4A_49_F8_00_00_00},
//{10_10_13_12_12_12_12_FF_12_12_12_12_13_10_10_00},/*"单",0*/
/* (16 X 16 , 宋体 )*/
			rdata_top<=128'h00_00_F8_49_4A_4C_48_F8_48_4C_4A_49_F8_00_00_00;
			rdata_btm<=128'h10_10_13_12_12_12_12_FF_12_12_12_12_13_10_10_00;
			end
		5'd1:begin
//{40_40_42_44_58_C0_40_7F_40_C0_50_48_46_40_40_00},
//{80_80_40_20_18_07_00_00_00_3F_40_40_40_40_78_00},/*"光",0*/
/* (16 X 16 , 宋体 )*/
			rdata_top<=128'h40_40_42_44_58_C0_40_7F_40_C0_50_48_46_40_40_00;
			rdata_btm<=128'h80_80_40_20_18_07_00_00_00_3F_40_40_40_40_78_00;
			end
		5'd2:begin
//{80_82_82_82_82_82_82_E2_A2_92_8A_86_82_80_80_00},
//{00_00_00_00_00_40_80_7F_00_00_00_00_00_00_00_00},/*"子",0*/
/* (16 X 16 , 宋体 )*/
			rdata_top<=128'h80_82_82_82_82_82_82_E2_A2_92_8A_86_82_80_80_00;
			rdata_btm<=128'h00_00_00_00_00_40_80_7F_00_00_00_00_00_00_00_00;
			end
		5'd3:begin
//{40_40_42_CC_00_40_40_40_40_FF_40_40_40_40_40_00},
//{00_00_00_7F_20_10_00_00_00_FF_00_00_00_00_00_00},/*"计",0*/
/* (16 X 16 , 宋体 )*/
			rdata_top<=128'h40_40_42_CC_00_40_40_40_40_FF_40_40_40_40_40_00;
			rdata_btm<=128'h00_00_00_7F_20_10_00_00_00_FF_00_00_00_00_00_00;
			end
		5'd4:begin
//{90_52_34_10_FF_10_34_52_80_70_8F_08_08_F8_08_00},
//{82_9A_56_63_22_52_8E_00_80_40_33_0C_33_40_80_00},/*"数",0*/
/* (16 X 16 , 宋体 )*/
			rdata_top<=128'h90_52_34_10_FF_10_34_52_80_70_8F_08_08_F8_08_00;
			rdata_btm<=128'h82_9A_56_63_22_52_8E_00_80_40_33_0C_33_40_80_00;
			end
		5'd5:begin
//{80_80_9E_92_92_92_9E_E0_80_9E_B2_D2_92_9E_80_00},
//{08_08_F4_94_92_92_F1_00_01_F2_92_94_94_F8_08_00},/*"器",0*/
/* (16 X 16 , 宋体 )*/
			rdata_top<=128'h80_80_9E_92_92_92_9E_E0_80_9E_B2_D2_92_9E_80_00;
			rdata_btm<=128'h08_08_F4_94_92_92_F1_00_01_F2_92_94_94_F8_08_00;
			end
		5'd6:begin
//{00_E0_10_08_08_10_E0_00_00_0F_10_20_20_10_0F_00},/*"0",0*/
/* (8 X 16 ,宋体 )*/
			rdata_top<=128'h00_E0_10_08_08_10_E0_00_00_00_00_00_00_00_00_00;
			rdata_btm<=128'h00_0F_10_20_20_10_0F_00_00_00_00_00_00_00_00_00;
			end
		5'd7:begin
//{00_00_10_10_F8_00_00_00_00_00_20_20_3F_20_20_00},/*"1",0*/
/* (8 X 16 , 宋体 )*/
			rdata_top<=128'h00_00_10_10_F8_00_00_00_00_00_00_00_00_00_00_00;
			rdata_btm<=128'h00_00_20_20_3F_20_20_00_00_00_00_00_00_00_00_00;
			end
		5'd8:begin
//{00_70_08_08_08_08_F0_00_00_30_28_24_22_21_30_00},/*"2",0*/
/* (8 X 16 , 宋体 )*/
			rdata_top<=128'h00_70_08_08_08_08_F0_00_00_00_00_00_00_00_00_00;
			rdata_btm<=128'h00_30_28_24_22_21_30_00_00_00_00_00_00_00_00_00;
			end
		5'd9:begin
//{00_30_08_08_08_88_70_00_00_18_20_21_21_22_1C_00},/*"3",0*/
/* (8 X 16 , 宋体 )*/
			rdata_top<=128'h00_30_08_08_08_88_70_00_00_00_00_00_00_00_00_00;
			rdata_btm<=128'h00_18_20_21_21_22_1C_00_00_00_00_00_00_00_00_00;
			end
		5'd10:begin
//{00_00_80_40_30_F8_00_00_00_06_05_24_24_3F_24_24},/*"4",0*/
/* (8 X 16 , 宋体 )*/
			rdata_top<=128'h00_00_80_40_30_F8_00_00_00_00_00_00_00_00_00_00;
			rdata_btm<=128'h00_06_05_24_24_3F_24_24_00_00_00_00_00_00_00_00;
			end
		5'd11:begin
//{00_F8_88_88_88_08_08_00_00_19_20_20_20_11_0E_00},/*"5",0*/
/* (8 X 16 , 宋体 )*/
			rdata_top<=128'h00_F8_88_88_88_08_08_00_00_00_00_00_00_00_00_00;
			rdata_btm<=128'h00_19_20_20_20_11_0E_00_00_00_00_00_00_00_00_00;
			end
		5'd12:begin
//{00_E0_10_88_88_90_00_00_00_0F_11_20_20_20_1F_00},/*"6",0*/
/* (8 X 16 , 宋体 )*/
			rdata_top<=128'h00_E0_10_88_88_90_00_00_00_00_00_00_00_00_00_00;
			rdata_btm<=128'h00_0F_11_20_20_20_1F_00_00_00_00_00_00_00_00_00;
			end
		5'd13:begin
//{00_18_08_08_88_68_18_00_00_00_00_3E_01_00_00_00},/*"7",0*/
/* (8 X 16 , 宋体 )*/
			rdata_top<=128'h00_18_08_08_88_68_18_00_00_00_00_00_00_00_00_00;
			rdata_btm<=128'h00_00_00_3E_01_00_00_00_00_00_00_00_00_00_00_00;
			end
		5'd14:begin
//{00_70_88_08_08_88_70_00_00_1C_22_21_21_22_1C_00},/*"8",0*/
/* (8 X 16 , 宋体 )*/
			rdata_top<=128'h00_70_88_08_08_88_70_00_00_00_00_00_00_00_00_00;
			rdata_btm<=128'h00_1C_22_21_21_22_1C_00_00_00_00_00_00_00_00_00;
			end
		5'd15:begin
//{00_F0_08_08_08_10_E0_00_00_01_12_22_22_11_0F_00},/*"9",0*/
/* (8 X 16 , 宋体 )*/
			rdata_top<=128'h00_F0_08_08_08_10_E0_00_00_00_00_00_00_00_00_00;
			rdata_btm<=128'h00_01_12_22_22_11_0F_00_00_00_00_00_00_00_00_00;
			end
		5'd16:begin
//{10_60_02_8C_00_44_54_54_54_7F_54_54_54_44_40_00}
//{04_04_7E_01_00_00_FF_15_15_15_55_95_7F_00_00_00}"清",0*/
/* (16 X 16 , 宋体 )*/
			rdata_top<=128'h10_60_02_8C_00_44_54_54_54_7F_54_54_54_44_40_00;
			rdata_btm<=128'h04_04_7E_01_00_00_FF_15_15_15_55_95_7F_00_00_00;
			end
		default:begin
					rdata_top<=128'd0;
					rdata_btm<=128'd0;
				end
	 endcase

assign data_top=rdata_top;
assign data_btm=rdata_btm;
endmodule
